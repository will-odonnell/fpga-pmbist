library verilog;
use verilog.vl_types.all;
entity mbist_top is
    generic(
        dw              : integer := 8;
        mw              : integer := 4;
        rw              : integer := 4;
        sw              : integer := 37;
        tasw            : integer := 8;
        tcsw            : integer := 4;
        tdsw            : integer := 8;
        spl_admd        : integer := 0;
        sph_admd        : integer := 3;
        spl_w           : integer := 4;
        sph_w           : integer := 4;
        spl_data        : integer := 5;
        sph_data        : integer := 12;
        spl_no          : integer := 13;
        sph_no          : integer := 14;
        spl_pol         : integer := 15;
        sph_pol         : integer := 18;
        spl_op          : integer := 19;
        sph_op          : integer := 34;
        spl_updwn       : integer := 35;
        sph_updwn       : integer := 35;
        sw_admd         : integer := 4;
        sw_w            : integer := 1;
        sw_data         : integer := 8;
        sw_no           : integer := 2;
        sw_pol          : integer := 4;
        sw_op           : integer := 16;
        sw_updwn        : integer := 1;
        irl_te          : integer := 0;
        irh_te          : integer := 0;
        irl_admd        : integer := 1;
        irh_admd        : integer := 4;
        irl_w           : integer := 5;
        irh_w           : integer := 5;
        irl_data        : integer := 6;
        irh_data        : integer := 13;
        irl_no          : integer := 14;
        irh_no          : integer := 15;
        irl_pol         : integer := 16;
        irh_pol         : integer := 19;
        irl_op          : integer := 20;
        irh_op          : integer := 35;
        irl_updwn       : integer := 36;
        irh_updwn       : integer := 36;
        irw_te          : integer := 1;
        irw_admd        : integer := 4;
        irw_w           : integer := 1;
        irw_data        : integer := 8;
        irw_no          : integer := 2;
        irw_pol         : integer := 4;
        irw_op          : integer := 16;
        irw_updwn       : integer := 1
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        ts_in           : in     vl_logic;
        scan_in         : in     vl_logic_vector;
        tas_out         : out    vl_logic_vector;
        tcs_out         : out    vl_logic_vector;
        tds_out         : out    vl_logic_vector;
        passfail_out    : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of dw : constant is 1;
    attribute mti_svvh_generic_type of mw : constant is 1;
    attribute mti_svvh_generic_type of rw : constant is 1;
    attribute mti_svvh_generic_type of sw : constant is 1;
    attribute mti_svvh_generic_type of tasw : constant is 1;
    attribute mti_svvh_generic_type of tcsw : constant is 1;
    attribute mti_svvh_generic_type of tdsw : constant is 1;
    attribute mti_svvh_generic_type of spl_admd : constant is 1;
    attribute mti_svvh_generic_type of sph_admd : constant is 1;
    attribute mti_svvh_generic_type of spl_w : constant is 1;
    attribute mti_svvh_generic_type of sph_w : constant is 1;
    attribute mti_svvh_generic_type of spl_data : constant is 1;
    attribute mti_svvh_generic_type of sph_data : constant is 1;
    attribute mti_svvh_generic_type of spl_no : constant is 1;
    attribute mti_svvh_generic_type of sph_no : constant is 1;
    attribute mti_svvh_generic_type of spl_pol : constant is 1;
    attribute mti_svvh_generic_type of sph_pol : constant is 1;
    attribute mti_svvh_generic_type of spl_op : constant is 1;
    attribute mti_svvh_generic_type of sph_op : constant is 1;
    attribute mti_svvh_generic_type of spl_updwn : constant is 1;
    attribute mti_svvh_generic_type of sph_updwn : constant is 1;
    attribute mti_svvh_generic_type of sw_admd : constant is 1;
    attribute mti_svvh_generic_type of sw_w : constant is 1;
    attribute mti_svvh_generic_type of sw_data : constant is 1;
    attribute mti_svvh_generic_type of sw_no : constant is 1;
    attribute mti_svvh_generic_type of sw_pol : constant is 1;
    attribute mti_svvh_generic_type of sw_op : constant is 1;
    attribute mti_svvh_generic_type of sw_updwn : constant is 1;
    attribute mti_svvh_generic_type of irl_te : constant is 1;
    attribute mti_svvh_generic_type of irh_te : constant is 1;
    attribute mti_svvh_generic_type of irl_admd : constant is 1;
    attribute mti_svvh_generic_type of irh_admd : constant is 1;
    attribute mti_svvh_generic_type of irl_w : constant is 1;
    attribute mti_svvh_generic_type of irh_w : constant is 1;
    attribute mti_svvh_generic_type of irl_data : constant is 1;
    attribute mti_svvh_generic_type of irh_data : constant is 1;
    attribute mti_svvh_generic_type of irl_no : constant is 1;
    attribute mti_svvh_generic_type of irh_no : constant is 1;
    attribute mti_svvh_generic_type of irl_pol : constant is 1;
    attribute mti_svvh_generic_type of irh_pol : constant is 1;
    attribute mti_svvh_generic_type of irl_op : constant is 1;
    attribute mti_svvh_generic_type of irh_op : constant is 1;
    attribute mti_svvh_generic_type of irl_updwn : constant is 1;
    attribute mti_svvh_generic_type of irh_updwn : constant is 1;
    attribute mti_svvh_generic_type of irw_te : constant is 1;
    attribute mti_svvh_generic_type of irw_admd : constant is 1;
    attribute mti_svvh_generic_type of irw_w : constant is 1;
    attribute mti_svvh_generic_type of irw_data : constant is 1;
    attribute mti_svvh_generic_type of irw_no : constant is 1;
    attribute mti_svvh_generic_type of irw_pol : constant is 1;
    attribute mti_svvh_generic_type of irw_op : constant is 1;
    attribute mti_svvh_generic_type of irw_updwn : constant is 1;
end mbist_top;
