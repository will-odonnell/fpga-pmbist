library verilog;
use verilog.vl_types.all;
entity cycle_controller is
    generic(
        mw              : integer := 4;
        cs              : integer := 2;
        irl_te          : integer := 0;
        irh_te          : integer := 0;
        irl_admd        : integer := 1;
        irh_admd        : integer := 4;
        irl_w           : integer := 5;
        irh_w           : integer := 5;
        irl_data        : integer := 6;
        irh_data        : integer := 13;
        irl_no          : integer := 14;
        irh_no          : integer := 15;
        irl_pol         : integer := 16;
        irh_pol         : integer := 19;
        irl_op          : integer := 20;
        irh_op          : integer := 35;
        irl_updwn       : integer := 36;
        irh_updwn       : integer := 36;
        irw_te          : integer := 1;
        irw_admd        : integer := 4;
        irw_w           : integer := 1;
        irw_data        : integer := 8;
        irw_no          : integer := 2;
        irw_pol         : integer := 4;
        irw_op          : integer := 16;
        irw_updwn       : integer := 1;
        ccw_pol         : integer := 1;
        ccw_op          : integer := 4
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        op_in           : in     vl_logic_vector;
        pol_in          : in     vl_logic_vector;
        no_in           : in     vl_logic_vector;
        ts_in           : in     vl_logic;
        op_out          : out    vl_logic_vector;
        pol_out         : out    vl_logic_vector;
        cc_cmp_out      : out    vl_logic;
        cc_cmpff_out    : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of mw : constant is 1;
    attribute mti_svvh_generic_type of cs : constant is 1;
    attribute mti_svvh_generic_type of irl_te : constant is 1;
    attribute mti_svvh_generic_type of irh_te : constant is 1;
    attribute mti_svvh_generic_type of irl_admd : constant is 1;
    attribute mti_svvh_generic_type of irh_admd : constant is 1;
    attribute mti_svvh_generic_type of irl_w : constant is 1;
    attribute mti_svvh_generic_type of irh_w : constant is 1;
    attribute mti_svvh_generic_type of irl_data : constant is 1;
    attribute mti_svvh_generic_type of irh_data : constant is 1;
    attribute mti_svvh_generic_type of irl_no : constant is 1;
    attribute mti_svvh_generic_type of irh_no : constant is 1;
    attribute mti_svvh_generic_type of irl_pol : constant is 1;
    attribute mti_svvh_generic_type of irh_pol : constant is 1;
    attribute mti_svvh_generic_type of irl_op : constant is 1;
    attribute mti_svvh_generic_type of irh_op : constant is 1;
    attribute mti_svvh_generic_type of irl_updwn : constant is 1;
    attribute mti_svvh_generic_type of irh_updwn : constant is 1;
    attribute mti_svvh_generic_type of irw_te : constant is 1;
    attribute mti_svvh_generic_type of irw_admd : constant is 1;
    attribute mti_svvh_generic_type of irw_w : constant is 1;
    attribute mti_svvh_generic_type of irw_data : constant is 1;
    attribute mti_svvh_generic_type of irw_no : constant is 1;
    attribute mti_svvh_generic_type of irw_pol : constant is 1;
    attribute mti_svvh_generic_type of irw_op : constant is 1;
    attribute mti_svvh_generic_type of irw_updwn : constant is 1;
    attribute mti_svvh_generic_type of ccw_pol : constant is 1;
    attribute mti_svvh_generic_type of ccw_op : constant is 1;
end cycle_controller;
