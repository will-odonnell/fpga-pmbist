library verilog;
use verilog.vl_types.all;
entity pmbist_test is
end pmbist_test;
