`include "defines.v"

//***********************************************
// Module Name 
//***********************************************
module decode_logic(tas_in,lu_out,ld_out);

//-----------------------------------------------
// Parameters and Definitions
//-----------------------------------------------
parameter   tasw        = `ADDR_WIDTH;


//-----------------------------------------------
// Input/Output Signals
//-----------------------------------------------
input    [tasw-1:0]	tas_in;
output    		lu_out;
output     		ld_out;

//-----------------------------------------------
// Internal Signals
//-----------------------------------------------
assign lu_out = tas_in[0];
assign ld_out = tas_in[0];

//***********************************************
// Module definition
//***********************************************

endmodule 
