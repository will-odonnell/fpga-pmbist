//***********************************************
// Module Name 
//***********************************************
module operation_formatting(op_in,op_out);
`include "defines.v"
//-----------------------------------------------
// Parameters and Definitions
//-----------------------------------------------
parameter    opw        = `IR_BFW_OP_SING;

//-----------------------------------------------
// Input/Output Signals
//-----------------------------------------------
input        [opw-1:0]  op_in;
output       [opw-1:0]  op_out;

//-----------------------------------------------
// Internal Signals
//-----------------------------------------------
assign op_out = op_in;

//***********************************************
// Module definition
//***********************************************

endmodule 
